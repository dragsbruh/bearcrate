module main

fn main() {
	println('Hugs! Beware its a Bear!')
}
